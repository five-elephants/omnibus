package Bus_tb;
	`include "bus_transactor.sv"
endpackage
